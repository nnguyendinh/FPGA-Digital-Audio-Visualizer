module audio_display_top(
		input rst, 
		input clk, 
      input clk_adc,
		input start,
		output reg hsync, 
		output reg vsync, 
		output reg [3:0] red, 
		output reg [3:0] green, 
		output reg [3:0] blue,
		output [9:0] leds
	);

    wire [17:0] s0;
    wire [17:0] s1;
    wire [17:0] s2;
    wire [17:0] s3;
    wire [17:0] s4;
    wire [17:0] s5;
    wire [17:0] s6;
    wire [17:0] s7;
    wire [17:0] s8;
    wire [17:0] s9;
    wire [17:0] s10;
    wire [17:0] s11;
    wire [17:0] s12;
    wire [17:0] s13;
    wire [17:0] s14;
    wire [17:0] s15;

    reg [17:0] b0 = 0;
    reg [17:0] b1 = 0;
    reg [17:0] b2 = 0;
    reg [17:0] b3 = 0;
    reg [17:0] b4 = 0;
    reg [17:0] b5 = 0;
    reg [17:0] b6 = 0;
    reg [17:0] b7 = 0;
    reg [17:0] b8 = 0;
    reg [17:0] b9 = 0;
    reg [17:0] b10 = 0;
    reg [17:0] b11 = 0;
    reg [17:0] b12 = 0;
    reg [17:0] b13 = 0;
    reg [17:0] b14 = 0;
    reg [17:0] b15 = 0;

    localparam IDLE = 0;
	localparam START = 1;
	localparam SAMPLING = 2;
	localparam FFT = 3;
    localparam DONE = 4;

	reg [2:0] state = IDLE;
	reg [2:0] state_d = IDLE;
	
	wire clk_25;
	wire clk_sampling;
    reg sampling_start = 0;
	 wire sampling_done;

	pll clk_generator(clk, clk_25);
	
	assign leds[9:2] = s0[9:2];
	assign leds[1] = start;
	assign leds[0] = clk_sampling;

    mic_sampler sampler(.clk_25(clk_25), .clk_adc(clk_adc), .start(1'b1), .done(sampling_done), .s0(s0), 
                        .s1(s1), .s2(s2), .s3(s3), .s4(s4), .s5(s5), .s6(s6), .s7(s7), .s8(s8), 
                        .s9(s9), .s10(s10), .s11(s11), .s12(s12), .s13(s13), .s14(s14), .s15(s15), .clk_sampling(clk_sampling));

	vga display(.vgaclk(clk_25), .rst(rst), .hsync(hsync), .vsync(vsync), .red(red), .green(green), .blue(blue), 
            .bar0(b0), .bar1(b1), .bar2(b2), .bar3(b3), .bar4(b4), .bar5(b5), .bar6(b6), .bar7(b7), .bar8(b8), 
            .bar9(b9), .bar10(b10), .bar11(b11), .bar12(b12), .bar13(b13), .bar14(b14), .bar15(b15));

	always @(posedge clk_25) begin
        state <= state_d;

        if (rst) begin
            sampling_start <= 0;
            state <= IDLE;
        end
        else if (state == IDLE) begin
            sampling_start <= 0;
        end
        else if (state == START) begin
            sampling_start <= 1;
        end
        else if (state == SAMPLING) begin
            sampling_start <= 0;
        end
        else if (state == FFT) begin
            sampling_start <= 0;
        end
        else if (state == DONE) begin
            sampling_start <= 0;
            b0 <= s0;
            b1 <= s1;
            b2 <= s2;
            b3 <= s3;
            b4 <= s4;
            b5 <= s5;
            b6 <= s6;
            b7 <= s7;
            b8 <= s8;
            b9 <= s9;
            b10 <= s10;
            b11 <= s11;
            b12 <= s12;
            b13 <= s13;
            b14 <= s14;
            b15 <= s15;
        end
    end

    always_comb begin

        case(state)
            IDLE: begin
                if (vsync) begin
                    state_d = START;
                end
                else begin
                    state_d = IDLE;
                end
            end
            START: begin
                state_d = SAMPLING;
            end
            SAMPLING: begin
                if (sampling_done) begin
                    state_d = DONE;
                end
                else    
                    state_d = SAMPLING;
            end
            // FFT state not included in this test
            FFT: begin
                state_d = IDLE;
            end
            DONE: begin
                if (vsync == 0) begin
                    state_d = IDLE;
                end
                else begin
                    state_d = DONE;
                end
            end
        endcase
    end

endmodule
